module usb_controller();


endmodule